LIBRARY IEEE;
USE ieee.std_logic_1164.all;

ENTITY NAND1 IS
    PORT (i0, i1: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	o: OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END ENTITY NAND1;

ARCHITECTURE Behavior OF NAND1 IS
    BEGIN
	outputs: FOR i IN 0 TO 31 GENERATE
     	    output: ENTITY work.NAND0(Behavior) PORT MAP (i0(i), i1(i), o(i));
	END GENERATE;
END ARCHITECTURE Behavior;
